module top(
	input clk,
	input rst
);
	datapath DP();
	controller CT();
endmodule