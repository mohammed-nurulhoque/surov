module controller();
endmodule 